// ALU codes for all possible ALU operations
// 4-bits wide
// Based off of the returned funct3/7 of the RISCV compiler
// https://riscvasm.lucasteske.dev/#
// both inputs will always be 32-bits
// input switching performed by decoder
// decoding immediates done via decoder switching

// ADD, code used for ADD and ADDI ins
// Adds two operands
`define ADD     4'd0

// SLT, set-less-than, used for STLI and STL
// result is 1 if operand1 < operand2 signed comparison, else 0
`define SLT     4'd2

// SLTU, set-less-than-unsigned, used for STLIU and STLU
// result is 1 if operand1 < operand2 unsigned comparison, else 0
`define SLTU    4'd3

// AND, logical and, used for AND and ANDI
// logically ANDs two operands together
`define AND     4'd7

// OR, logical or, used for OR and ORI
// logically ORs two operands together
`define OR      4'd6

// XOR, logical xor, used for XOR and XORI
// logically XORs two operands together
`define XOR     4'd4

// SLL, shift-left-logical, used for SLL and SLLI
// logically shifts first operand left by second
// (zeros shifted into lower bits)
// Will only use lower 5 bits of second operand
`define SLL     4'd1

// SRL, shift-right-logical, used for SRL and SRLI
// logically shifts first operand right by second
// (zeros shifted into upper bits)
// Will only use lower 5 bits of second operand
`define SRL     4'd5

// SRA, shift-right-arithemetic, used for SRA and SRAI
// arithemetically shifts first operand right by second
// (sign bit is shifted into upper bits)
// Will only use lower 5 bits of second operand
`define SRA     4'd13
// NOTE: on immediate opcode, shares a funct3 with SRL, system will include rawIns[30] as MSB of opcode

// SUB, subtract, used for SUB
// subtracts the first operand from the second
// only exists as an R-type instruction
`define SUB     4'd8

// CPY, repeats the value in operand 2, used for LUI
`define CPY     4'b1111