// Instruction codes for constant zero argument instructions
`define NOP 32'b0000_0000_0000_0000_0000_0000_0000_0011