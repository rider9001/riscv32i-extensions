// Multplication codes file

`define MULC     2'd0

`define MULHC    2'd1

`define MULHUC   2'd2

`define MULHSUC  2'd3