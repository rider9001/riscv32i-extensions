// Division codes file

`define DIVC    2'd0

`define REMC    2'd1

`define DIVUC   2'd2

`define REMUC   2'd3