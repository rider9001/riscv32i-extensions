// Zero delay RAM module
// implemented as a test tool for the RSICV32I processor
// Will try implementing a multi-cycle RAM later
// Takes the address of the LSBtye and returns 4 bytes
// Stores all data as bytes, any read lower than 4 is invalid
// First 16 bytes are reserved as hardware async input/output addresses
// 0x0 = Inp1, 0x4 = Inp2, 0x8 = Out1, 0xB = Out2
module zeroDelayRAM #(parameter dataW = 32, parameter RAMAddrSize = 32)
(
    input logic clock, reset,
    input logic [RAMAddrSize-1:0] RAMAddr,
    input logic [dataW-1:0] DataIn,
    input logic WriteControl,
    input logic [dataW-1:0] UsrInpData1, UsrInpData2,
    output logic [dataW-1:0] DataOut,
    output logic [dataW-1:0] UsrOutData1, UsrOutData2
);

timeunit 1ns; timeprecision 10ps;

// Create version of RAM address shifted into 4 byte per-unit range
logic [RAMAddrSize-1:0] RAMAddrAdj;
assign RAMAddrAdj = RAMAddr>>2;

logic [dataW-1:0] RAMArray [3:(1<<(RAMAddrSize>>2))];

always_comb
begin
    case (RAMAddrAdj)
        0: DataOut = UsrInpData1;
        1: DataOut = UsrInpData2;
        2: DataOut = UsrOutData1;
        3: DataOut = UsrOutData2;
        default: DataOut = RAMArray[RAMAddrAdj];
    endcase
end

always_ff @( posedge clock, posedge reset )
begin
    if (reset)  RAMArray <= '{default: '0};
    else
    begin
        // Writes to input sectors are blocked
        if (WriteControl && RAMAddrAdj > 1)
        begin
            case (RAMAddrAdj)
                2: UsrOutData1 <= DataIn;
                3: UsrOutData2 <= DataIn;
                default: RAMArray[RAMAddrAdj] <= DataIn;
            endcase
        end
    end
end

endmodule